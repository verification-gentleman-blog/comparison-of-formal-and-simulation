// Copyright 2020 Tudor Timisescu (verificationgentleman.com)
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.


class reserved_ctrl_values_coverage;

  covergroup cg with function sample(bit [1:0] shape, bit [5:0] operation);
    coverpoint shape {
      ignore_bins keep = { RECTANGLE, TRIANGLE, KEEP_SHAPE };
    }
    coverpoint operation {
      ignore_bins keep = {
          PERIMETER, AREA, IS_SQUARE, IS_EQUILATERAL, IS_ISOSCELES, KEEP_OPERATION };
    }
  endgroup


  function new();
    cg = new();
  endfunction


  function void sample(uvm_reg_data_t SHAPE, uvm_reg_data_t OPERATION);
    cg.sample(SHAPE, OPERATION);
  endfunction

endclass
