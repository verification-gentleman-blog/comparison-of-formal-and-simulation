// Copyright 2020 Tudor Timisescu (verificationgentleman.com)
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.


package shape_processor_tests;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "reg_access_macros.svh"

  `include "virtual_sequencer.svh"
  `include "abstract_test.svh"

  `include "random_ctrl_writes.svh"
  `include "random_ctrl_writes_with_nonreserved_values.svh"
  `include "random_ctrl_writes_with_reserved_shape_values.svh"
  `include "random_ctrl_writes_with_reserved_operation_values.svh"

endpackage
