// Copyright 2020 Tudor Timisescu (verificationgentleman.com)
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.


module shape_processor_props(
    input bit rst_n,
    input bit clk,

    input bit write,
    input bit [31:0] write_data,

    input bit read,
    input bit [31:0] read_data,

    input bit error,

    input bit [31:0] ctrl_sfr
    );

  default disable iff !rst_n;

  default clocking @(posedge clk);
  endclocking


  write_data_written_to_ctrl_sfr: assert property (
      write |=> ctrl_sfr == $past(write_data)
      );

  ctrl_sfr_constant_if_no_write: assert property (
      !write |=> $stable(ctrl_sfr)
      );

endmodule


bind shape_processor shape_processor_props props(.*);
