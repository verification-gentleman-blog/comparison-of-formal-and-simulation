// Copyright 2020 Tudor Timisescu (verificationgentleman.com)
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.


`include "coverage/ctrl_value_combinations_coverage.svh"
`include "coverage/legal_ctrl_value_combinations_coverage.svh"
`include "coverage/illegal_ctrl_value_combinations_coverage.svh"
`include "coverage/reserved_ctrl_values_coverage.svh"
`include "coverage/ctrl_coverage_collector.svh"

`include "coverage/ctrl_keep_operation_value_combinations_coverage.svh"
`include "coverage/ctrl_keep_operation_coverage_collector.svh"

`include "coverage/ctrl_keep_both_coverage_collector.svh"
