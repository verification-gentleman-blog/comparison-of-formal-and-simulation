// Copyright 2020 Tudor Timisescu (verificationgentleman.com)
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.


class test_ctrl_sequence extends uvm_sequence;

  function new(string name = get_type_name());
    super.new(name);
  endfunction


  virtual task body();
    write_ctrl_values_sequence write_ctrl_values;
    `uvm_do(write_ctrl_values)
    `read_reg(p_sequencer.regs.CTRL)
  endtask


  `uvm_object_utils(test_ctrl_sequence)
  `uvm_declare_p_sequencer(virtual_sequencer)

endclass
